`timescale 1ns/1ns

module tb; //testbench module

integer input_file, output_file, in, out;
integer i;

parameter CYCLE = 100;

reg clk, reset_n;
reg start, done;
reg [31:0] a_in, b_in;
reg [31:0] result;


//clock generation for write clock
initial begin
  clk <= 0;
  forever #(CYCLE/2) clk = ~clk;
end

//release of reset_n relative to two clocks
initial begin
    input_file  = $fopen("input_data", "rb");
    if (input_file==0) begin
      $display("ERROR : CAN NOT OPEN input_file");
    end
    output_file = $fopen("output_data", "wb");
    if (output_file==0) begin
      $display("ERROR : CAN NOT OPEN output_file");
    end
    a_in='x;
    b_in='x;
    start=1'b0;
    reset_n <= 0;
    #(CYCLE * 1.5) reset_n = 1'b1; //reset for 1.5 clock cycles
end

gcd gcd_0(.*); //instantiate the gcd unit

initial begin

  #(CYCLE*4);  //delay after reset
  while(! $feof(input_file)) begin
   $fscanf(input_file,"%d %d", a_in, b_in);
   start=1'b1;
   #(CYCLE);
   start=1'b0;
   while(done != 1'b1) #(CYCLE);
   $display ("a_in=%d   b_in=%d   result=%d", a_in, b_in, result);
   $fwrite(output_file,"a_in	b_in	result\n");
   $fwrite(output_file,"%d	%d	%d\n",a_in,b_in, result);
   #(CYCLE*2); //2 cycle delay between trials
  end
$stop;
$fclose(input_file);
end

endmodule
